module CUMULATIVE_ADDER(
	DATA_IN,
	DATA_OUT,
	TRIGGER
);

/*

DATA_IN 14 bits

*/

input DATA_IN;
output DATA_OUT;
output TRIGGER;